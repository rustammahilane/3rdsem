module not_(
	input a,
	output y
);
assign y = ~a;
endmodule
